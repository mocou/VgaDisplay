module VgaDisplay(
			clk,
			rst,
			en
		);


endmodule
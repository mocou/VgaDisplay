module VgaDisplay(
			
		);


endmodule